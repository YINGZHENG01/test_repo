module key
(


);



endmodule
